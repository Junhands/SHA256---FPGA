`default_nettype none
module CLA_cell(
    input  wire a,
    input  wire b,
    input  wire c_in,
    output wire c_out,
    output wire sum
);
    